module hello_ModuleA;
    initial begin
        $display("Hello, world!");
    end
endmodule
